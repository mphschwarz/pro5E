// SPI Treiber für die IO-Expander MCP23S17
// \_toolchain\datasheets\MCP23S17.pdf
module CLIENT_MCP23S17(
	input CLK,
	input SPI_MISO,
	input [15:0] IO16_D,
	output wire SPI_CS,
	output wire SPI_CLK,
	output wire SPI_MOSI,
	output reg [15:0] IO16_SW
	);
	//
	// Registerdefinition MCP23S17
	localparam IODIRA    = 8'h00; //Data Direction Register for PORTA   
	localparam IODIRB    = 8'h01; //Data Direction Register for PORTB
	localparam IPOLA     = 8'h02; //Input Polarity Register for PORTA
	localparam IPOLB     = 8'h03; //Input Polarity Register for PORTB
	localparam GPINTENA  = 8'h04; //Interrupt-on-change enable Register for PORTA
	localparam GPINTENB  = 8'h05; //Interrupt-on-change enable Register for PORTB
	localparam DEFVALA   = 8'h06; //Default Value Register for PORTA   
	localparam DEFVALB   = 8'h07; //Default Value Register for PORTB     
	localparam INTCONA   = 8'h08; //Interrupt-on-change control Register for PORTA 
	localparam INTCONB   = 8'h09; //Interrupt-on-change control Register for PORTB     
	localparam IOCON     = 8'h0A; //Configuration register for device                     
	localparam GPPUA     = 8'h0C; //100kOhm pullup resistor register for PORTA (sets pin to input when set)   
	localparam GPPUB     = 8'h0D; //100kOhm pullup resistor register for PORTB (sets pin to input when set)     
	localparam INTFA     = 8'h0E; //Interrupt flag Register for PORTA       
	localparam INTFB     = 8'h0F; //Interrupt flag Register for PORTB   
	localparam INTCAPA   = 8'h10; //Interrupt captured value Register for PORTA 
	localparam INTCAPB   = 8'h11; //Interrupt captured value Register for PORTB   
	localparam GPIOA     = 8'h12; //General purpose I/O Register for PORTA 
	localparam GPIOB     = 8'h13; //General purpose I/O Register for PORTB
	localparam OLATA     = 8'h14; //Output latch Register for PORTA
	localparam OLATB     = 8'h15; //Output latch Register for PORTB  	
	//
	// Read Write U1 und U2
	localparam R_U1 = 8'h4B;// 0x4B Adresse 5
	localparam W_U1 = 8'h4A;// 0x4A Adresse 5
	localparam R_U2 = 8'h4D;// 0x4D Adresse 6
	localparam W_U2 = 8'h4C;// 0x4C Adresse 6 
	//
	//localparam INIT = 3'd0;
	//
	reg [4:0] state;
	reg start;
	wire [23:0] data_in;
	reg [23:0] data_out;
	reg [15:0] counter;
	wire done;
	reg hri1; reg hri2; reg hri3; reg hri4; reg hri5; reg hri6;
	wire done_re; wire done_fe;
	//
	assign done_re = (hri1 && !hri2);
	assign done_fe = (!hri1 && hri2);
	//
	SPI_INP_FILTER_CLIENT spi_inp_filter_miso(CLK, SPI_MISO, spi_miso_filter); 
	defparam spi_inp_filter_miso.FILTER = 5'd2;
	SHIFTER_24_BIT shifter_24_bit(CLK, start, spi_miso_filter, data_out, done, SPI_CS, SPI_CLK, SPI_MOSI, data_in); 
	defparam shifter_24_bit.CLK_COUNTER = 5'd50;// 500kHz
	//
	initial
	begin
		//
		counter <= 0;
		state <= 0;
		data_out <= 0;
		start <= 0;
		hri1 <= 0; hri2 <= 0; hri3 <= 0; hri4 <= 0; hri5 <= 0; hri6 <= 0;
	end
	//
	
	//
	always @(posedge CLK)
	begin
	//
	hri1 <= done;
	hri2 <= hri1;
	//
	if (state == 0)
		begin
		start <= 0;
		state <= state + 1;
		end
	//
	if (state == 1)
		begin
		counter <= counter + 1;
		if (counter > 1000)
			begin
			counter <= 0;
			state <= state + 1;
			end
		end
	//
	if (state == 2) /* sequential operation mode disabled, address mode enabled */
	begin
		data_out[23:16] <= 8'h40; data_out[15:08] <= IOCON;	data_out[07:00] <= 8'h28;
		start <= 1;
		if (done_re) state <= state + 1;
	end
	//
	if (state == 3) begin start <= 0; state <= state + 1; end
	//
	if (state == 4) /* sequential operation mode disabled, address mode enabled */
	begin
		data_out[23:16] <= W_U1; data_out[15:08] <= IOCON;	data_out[07:00] <= 8'h28;
		start <= 1;
		if (done_re) state <= state + 1;
	end
	//
	if (state == 5) begin start <= 0; state <= state + 1; end
	//
	if (state == 6) /* sequential operation mode disabled, address mode enabled */
	begin
		data_out[23:16] <= W_U2; data_out[15:08] <= IOCON;	data_out[07:00] <= 8'h28;
		start <= 1;
		if (done_re) state <= state + 1;
	end
	//
	if (state == 7) begin start <= 0; state <= state + 1; end
	//
	if (state == 8) /* 1 = GPIO register bit will reflect the opposite logic state of the input pin. 0 = GPIO register bit will reflect the same logic state of the input pin. */
	begin
		data_out[23:16] <= W_U1; data_out[15:08] <= IPOLA;	data_out[07:00] <= 8'hFF;
		start <= 1;
		if (done_re) state <= state + 1;
	end
	//
	if (state == 9) begin start <= 0; state <= state + 1; end
	//
	if (state == 10) /* 1 = GPIO register bit will reflect the opposite logic state of the input pin. 0 = GPIO register bit will reflect the same logic state of the input pin. */
	begin
		data_out[23:16] <= W_U2; data_out[15:08] <= IPOLA;	data_out[07:00] <= 8'hFF;
		start <= 1;
		if (done_re) state <= state + 1;
	end
	//
	if (state == 11) begin start <= 0; state <= state + 1; end
	//
	if (state == 12) /* direction PORT A, 0 = OUTPUT, 1 = INPUT */
	begin
		data_out[23:16] <= W_U1; data_out[15:08] <= IODIRA;	data_out[07:00] <= 8'hFF;
		start <= 1;
		if (done_re) state <= state + 1;
	end
	//
	if (state == 13) begin start <= 0; state <= state + 1; end
	//
	if (state == 14) /* direction PORT B, 0 = OUTPUT, 1 = INPUT */
	begin
		data_out[23:16] <= W_U1; data_out[15:08] <= IODIRB;	data_out[07:00] <= 8'h00;
		start <= 1;
		if (done_re) state <= state + 1;
	end
	//
	if (state == 15) begin start <= 0; state <= state + 1; end
	//
	if (state == 16) /* direction PORT A, 0 = OUTPUT, 1 = INPUT */
	begin
		data_out[23:16] <= W_U2; data_out[15:08] <= IODIRA;	data_out[07:00] <= 8'hFF;
		start <= 1;
		if (done_re) state <= state + 1;
	end
	//
	if (state == 17) begin start <= 0; state <= state + 1; end
	//
	if (state == 18) /* direction PORT B, 0 = OUTPUT, 1 = INPUT */
	begin
		data_out[23:16] <= W_U2; data_out[15:08] <= IODIRB;	data_out[07:00] <= 8'h00;
		start <= 1;
		if (done_re) state <= state + 1;
	end
	//
	////////////////////////////////////////////////	
	if (state == 19) begin start <= 0; state <= state + 1; end
	//
	if (state == 20) /* read INPUTS */
	begin
		data_out[23:16] <= R_U1; data_out[15:08] <= GPIOA;	data_out[07:00] <= 8'hFF;
		IO16_SW[7:0] <= data_in[07:00];
		start <= 1;
		if (done_re) state <= state + 1;
	end
	//
	if (state == 21) begin start <= 0; state <= state + 1; end
	//
	if (state == 22) /* write OUTPUTS */
	begin
		data_out[23:16] <= W_U1; data_out[15:08] <= GPIOB;	data_out[07:00] <= IO16_D[7:0];
		start <= 1;
		if (done_re) state <= state + 1;
	end
	////////////////////////////////////////////////	
	if (state == 23) begin start <= 0; state <= state + 1; end
	//
	if (state == 24) /* read INPUTS */
	begin
		data_out[23:16] <= R_U2; data_out[15:08] <= GPIOA;	data_out[07:00] <= 8'hFF;
		IO16_SW[15:8] <= data_in[07:00];
		start <= 1;
		if (done_re) state <= state + 1;
	end
	//	
	if (state == 25) begin start <= 0; state <= state + 1; end
	//
	if (state == 26) /* write OUTPUTS */
	begin
		data_out[23:16] <= W_U2; data_out[15:08] <= GPIOB;	data_out[07:00] <= IO16_D[15:8];
		start <= 1;
		if (done_re) state <= 19;
	end
	////////////////////////////////////////////////		
	end
endmodule
////////////////////////////////////////////////////////////////////////////////////////////
//	24-BIT-Shifter
module SHIFTER_24_BIT(
	input CLK,
	input START,
	input IO_IN,
	input [23:0] DATA_OUT,
	output reg DONE,
	output reg CS,
	output reg CLK_OUT,
	output reg IO_OUT,
	output reg [23:0] DATA_IN
	);
	//
	parameter CLK_COUNTER = 5'd25;// 1MHz
	//
	reg [7:0] state;
	reg	[15:0]counter;
	reg	[15:0]counter_cs;
	reg enable;
	reg [7:0] clk_counter;
	reg [7:0] in_counter;
	reg [7:0] out_counter;	
	reg hri1; reg hri2; reg hri3; reg hri4;
	wire start_re; wire start_fe;
	wire clk_out_re; wire clk_out_fe;
	//
	assign start_re = (hri1 && !hri2);
	assign start_fe = (!hri1 && hri2);
	assign clk_out_re = (hri3 && !hri4);
	assign clk_out_fe = (!hri3 && hri4);	
	//
	initial
	begin
		DONE <= 0;
		CS <= 1;
		CLK_OUT <= 0;
		IO_OUT <= 0;
		DATA_IN <= 0;
		//
		state <= 0;
		counter <= 0;
		enable <= 0;
		clk_counter <= 0;
		in_counter <= 23;
		out_counter <= 23;
		counter_cs <= 0;
		hri1 <= 0; hri2 <= 0; hri3 <= 0; hri4 <= 0;
	end
	//
	always @(posedge CLK)
	begin
	//
	hri1 <= START;
	hri2 <= hri1;
	hri3 <= CLK_OUT;
	hri4 <= hri3;	
	//
	if (state == 0)
		begin
		counter_cs <= 0;
		clk_counter <= 0;
		in_counter <= 23;
		out_counter <= 23;
		if (start_re) 
			begin
			CS <= 0;
			DONE <= 0;
			state <= state + 1;		
			end
		//
		end
	//
	if (state == 1)
		begin
		counter_cs <= counter_cs + 1;
		if (counter_cs > 100) 
			begin
			counter_cs <= 0;
			enable <= 1;
			state <= state + 1;		
			end
		//
		end
	//
	if (state == 2)
		begin
		if (clk_counter == 48) 
			begin
			enable <= 0;
			state <= state + 1;		
			end
		//
		end
	//
	if (state == 3)
		begin
		counter_cs <= counter_cs + 1;
		if (counter_cs > 100) 
			begin
			counter_cs <= 0;
			CS <= 1;
			state <= state + 1;		
			end
		//
		end
	//
	if (state == 4)
		begin
		counter_cs <= counter_cs + 1;
		if (counter_cs > 100) 
			begin
			counter_cs <= 0;
			DONE <= 1;
			state <= 0;		
			end
		//
		end
	//
	////////////////////////////////////////////
	if (clk_out_re)
		begin
		DATA_IN[in_counter] <= IO_IN;
		if (in_counter > 0) in_counter <= in_counter - 1;
		end
	////////////////////////////////////////////
	IO_OUT <= DATA_OUT[out_counter];
	if (clk_out_fe)
		begin
		if (out_counter > 0) out_counter <= out_counter - 1;
		end
	////////////////////////////////////////////
	// Clockgenerator
	if (enable) 
		begin
		counter <= counter + 1;
		if(enable && (counter == CLK_COUNTER)) 
			begin
			counter <= 1;
			CLK_OUT <= !CLK_OUT;
			clk_counter <= clk_counter + 1;
			end	
		end
	else counter <= 1;
	//
	end
endmodule

////////////////////////////////////////////////////////////////////////////////////////////
//	Digitales Filter der Eingangssignale
module	SPI_INP_FILTER_CLIENT (
	input CLK, 
	input IN,
	output reg OUT
	);
//
parameter FILTER = 5'd10;
//
reg [4:0] ctr0;
reg [4:0] ctr1;
//
initial
	begin
	OUT <= 0;
	ctr0 <= 0;
	ctr1 <= 0;
	end
always	@(posedge CLK)
begin
	if (IN && !OUT)
		begin
		ctr0 <= 0;
		ctr1 <= ctr1 + 1;
		end
	//	
	if (!IN && OUT)
		begin
		ctr0 <= ctr0 + 1;
		ctr1 <= 0;
		end	
	//
	if (ctr0 == FILTER)
		begin
		ctr0 <= 0;
		ctr1 <= 0;
		OUT <= 0;
		end
	//
	if (ctr1 == FILTER)
		begin
		ctr0 <= 0;
		ctr1 <= 0;
		OUT <= 1;
		end
	//	
	if (((ctr0 > 0) && IN) || ((ctr1 > 0) && !IN))
		begin
		ctr0 <= 0;
		ctr1 <= 0;
		end	
end
endmodule
////////////////////////////////////////////////////////////////////////////////////////////
/*
ToDo: 
- FSM mit case
- Erweiterung PCB Tresor
- Beachtung der Warnungen bezüglich Datenbreite
- Signalfilter für die Eingangssignale der Tasten
*/
